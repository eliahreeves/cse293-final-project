// Implements CRC32 calculation for Ethernet FCS
// Used by packet_gen to add frame check sequences