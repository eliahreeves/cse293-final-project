// top module
// connects RMII (Reduced Media Independent Interface) to AXI Stream
// Instantiates packet_tx and packet_rx
