// Generates Ethernet/IP/UDP headers based on configured parameters
// Used by packet_gen to create valid network packets